module przesuniecie (
    ports
);
    
endmodule