//moduł porównania wartości sygnałów wejściowych A i B

module porownanie (i_arg_A, i_arg_B, o_result);
    parameter BITS = 32;
    
endmodule